/*
Description
Author : Foez Ahmed (foez.official@gmail.com)
*/

module rv_g_regfile_tb;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int XLEN = 64;
  localparam int FLEN = 32;
  localparam int MaxLen = (XLEN > FLEN) ? XLEN : FLEN;
  localparam bit AllowForwarding = 1;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns

  `CREATE_CLK(clk_i, 4ns, 6ns)
  logic              arst_ni = 1;
  logic [       5:0] wr_addr_i = '0;
  logic [MaxLen-1:0] wr_data_i = '0;
  logic              wr_en_i = '0;
  logic [       5:0] rd_addr_i = '0;
  logic [       5:0] rs1_addr_i = '0;
  logic [       5:0] rs2_addr_i = '0;
  logic [       5:0] rs3_addr_i = '0;
  logic              req_i = '0;
  logic [MaxLen-1:0] rs1_data_o;
  logic [MaxLen-1:0] rs2_data_o;
  logic [MaxLen-1:0] rs3_data_o;
  logic              gnt_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  rv_g_regfile #(
      .XLEN(XLEN),
      .FLEN(FLEN),
      .ALLOW_FORWARDING(AllowForwarding)
  ) u_rv_g_regfile (
      .arst_ni,
      .clk_i,
      .wr_addr_i,
      .wr_data_i,
      .wr_en_i,
      .rd_addr_i,
      .rs1_addr_i,
      .rs2_addr_i,
      .rs3_addr_i,
      .req_i,
      .rs1_data_o,
      .rs2_data_o,
      .rs3_data_o,
      .gnt_o
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100ns;
    arst_ni <= 0;
    #100ns;
    arst_ni <= 1;
    #100ns;
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    apply_reset();
    start_clk_i();

    @(posedge clk_i);
    result_print(1, "This is a Forced PASS");
    @(posedge clk_i);

    $finish;

  end

endmodule
