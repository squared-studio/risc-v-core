/*
Write a markdown documentation for this systemverilog module:
Author : Foez Ahmed (foez.official@gmail.com)
*/
`ifndef RV_G_PKG_SV__
`define RV_G_PKG_SV__

package rv_g_pkg;

  // NO IMMEDIATE
  `define NONE 3'b000

  // BTYPE INSTRUCTION IMMEDIATE
  `define BIMM 3'b001

  // ITYPE INSTRUCTION IMMEDIATE
  `define IIMM 3'b010

  // JTYPE INSTRUCTION IMMEDIATE
  `define JIMM 3'b011

  // RTYPE INSTRUCTION IMMEDIATE
  `define SIMM 3'b100

  // UTYPE INSTRUCTION IMMEDIATE
  `define UIMM 3'b101

  // CSR INSTRUCTION IMMEDIATE
  `define CIMM 3'b110

  `define _YES_ 1'b1
  `define _____ 1'b0

`ifdef READY__________________
  typedef enum logic [19:0] {
    //           EXTRA__  IMM__  frs3__  frs2__  frs1__  frd___  xrs2__  xrs1__  xrd___
    INVALID   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____},
    LUI       = {8'b0000_0000, `UIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_YES_},
    AUIPC     = {8'b0000_0000, `UIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_YES_},
    JAL       = {8'b0000_0000, `JIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_YES_},
    JALR      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    BEQ       = {8'b0000_0000, `BIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    BNE       = {8'b0000_0000, `BIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    BLT       = {8'b0000_0000, `BIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    BGE       = {8'b0000_0000, `BIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    BLTU      = {8'b0000_0000, `BIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    BGEU      = {8'b0000_0000, `BIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    LB        = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    LH        = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    LW        = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    LBU       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    LHU       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SB        = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    SH        = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    SW        = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    ADDI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SLTI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SLTIU     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    XORI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    ORI       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    ANDI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SLLI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SRLI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SRAI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    ADD       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SUB       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SLL       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SLT       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SLTU      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    XOR       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SRL       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SRA       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    OR        = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AND       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    FENCE     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    FENCE_TSO = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____},
    PAUSE     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____},
    ECALL     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____},
    EBREAK    = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____},
    LWU       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    LD        = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SD        = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_____},
    SLLI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SRLI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SRAI      = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    ADDIW     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SLLIW     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SRLIW     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SRAIW     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    ADDW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SUBW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SLLW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SRLW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    SRAW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    FENC_I    = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    CSRRW     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    CSRRS     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    CSRRC     = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    CSRRWI    = {8'b0000_0000, `CIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_YES_},
    CSRRSI    = {8'b0000_0000, `CIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_YES_},
    CSRRCI    = {8'b0000_0000, `CIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_YES_},
    MUL       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    MULH      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    MULHSU    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    MULHU     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    DIV       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    DIVU      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    REM       = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    REMU      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    MULW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    DIVW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    DIVUW     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    REMW      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    REMUW     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    LR_W      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SC_W      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOSWAP_W = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOADD_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOXOR_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOAND_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOOR_W   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMIN_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMAX_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMINU_W = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMAXU_W = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    LR_D      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    SC_D      = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOSWAP_D = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOADD_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOXOR_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOAND_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOOR_D   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMIN_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMAX_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMINU_D = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},
    AMOMAXU_D = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_YES_, `_YES_, `_YES_},

    FLW       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSW       = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMADD_S   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMSUB_S   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMSUB_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMADD_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FADD_S    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSUB_S    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMUL_S    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FDIV_S    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSQRT_S   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJ_S   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJN_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJX_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMIN_S    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMAX_S    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_W_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_WU_S = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMV_X_W   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FEQ_S     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLT_S     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLE_S     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCLASS_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_S_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_S_WU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMV_W_X   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_L_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_LU_S = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_S_L  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_S_LU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--

    FLD       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSD       = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMADD_D   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMSUB_D   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMSUB_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMADD_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FADD_D    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSUB_D    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMUL_D    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FDIV_D    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSQRT_D   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJ_D   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJN_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJX_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMIN_D    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMAX_D    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_S_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_D_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FEQ_D     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLT_D     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLE_D     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCLASS_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_W_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_WU_D = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_D_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_D_WU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_L_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_LU_D = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMV_X_D   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_D_L  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_D_LU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMV_D_X   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--

    FLQ       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSQ       = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMADD_Q   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMSUB_Q   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMSUB_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMADD_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FADD_Q    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSUB_Q    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMUL_Q    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FDIV_Q    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSQRT_Q   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJ_Q   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJN_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJX_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMIN_Q    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMAX_Q    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_S_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_Q_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_D_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_Q_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FEQ_Q     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLT_Q     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLE_Q     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCLASS_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_W_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_WU_Q = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_Q_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_Q_WU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_L_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_LU_Q = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_Q_L  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_Q_LU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--

    FLH       = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSH       = {8'b0000_0000, `SIMM, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMADD_H   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMSUB_H   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMSUB_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FNMADD_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FADD_H    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSUB_H    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMUL_H    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FDIV_H    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSQRT_H   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJ_H   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJN_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FSGNJX_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMIN_H    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMAX_H    = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_S_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_H_S  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_D_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_H_D  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_Q_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_H_Q  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FEQ_H     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLT_H     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FLE_H     = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCLASS_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_W_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_WU_H = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMV_X_H   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_H_W  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_H_WU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FMV_H_X   = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_L_H  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_LU_H = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_H_L  = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--
    FCVT_H_LU = {8'b0000_0000, `NONE, `_____, `_____, `_____, `_____, `_____, `_____, `_____}, //--

    WRS_NTO   = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_},
    WRS_STO   = {8'b0000_0000, `IIMM, `_____, `_____, `_____, `_____, `_____, `_YES_, `_YES_}
  } funct_t;
`endif

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

endpackage

`endif
