module tb_func_decode;
  initial begin
    $display("Hello!!");
  end
endmodule
